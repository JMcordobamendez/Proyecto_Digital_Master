library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Prueba integración de todo el Hardware junto :)
entity HARDWARE_1 is
    port(     CLK : in std_logic;
	        RESET : in std_logic;
			   RX : in std_logic;
		    HSYNC : out std_logic;
		    VSYNC : out std_logic;
	      COLOR_R : out std_logic_vector(3 downto 0);
	      COLOR_G : out std_logic_vector(3 downto 0);
	      COLOR_B : out std_logic_vector(3 downto 0));
end HARDWARE_1;
architecture A1 of HARDWARE_1 is
    --Define the components
    --Data path of the VGA
    component VGA_DATA is
	    port(    CLK : in std_logic;
	           DOUTB : in std_logic_vector(7 downto 0);
		       RESET : in std_logic;
		          CH : in std_logic_vector(9 downto 0);
		          CV : in std_logic_vector(9 downto 0);
		        ADDB : out std_logic_vector(9 downto 0);
		         ENB : out std_logic;
		       COLOR : out std_logic_vector(3 downto 0));
	end component;
	--Synchronizer/Controller of VGA
	component CONTROL_VGA is
	    port(    CLK : in std_logic;
	           RESET : in std_logic;
			   HSYNC : out std_logic;
			   VSYNC : out std_logic;
			    CH_o : out std_logic_vector(9 downto 0);
			    CV_o : out std_logic_vector(9 downto 0));
	end component;
	--Driver to read UART protocol
    component UART_RX is
    generic (
      BAUDRATE : INTEGER := 115200;     -- Desired baudrate
      CLK_FREQ : INTEGER := 100000000  -- Input clock in Hz
    );
    port (
      reset    : IN  STD_LOGIC;
      clk      : IN  STD_LOGIC;
      rx       : IN  STD_LOGIC;
      data_out : OUT STD_LOGIC_VECTOR (7 DOWNTO 0 );
      ready    : OUT STD_LOGIC
    );
    end component;
    --Driver to store the data of the UART in the RAM
    component CONTROL_UART is
    port( READY : in std_logic;
	      RESET : in std_logic;
		    CLK : in std_logic;
		   DATA : in std_logic_vector(7 downto 0);
		   ADDA : out std_logic_vector(9 downto 0);
		  ENA_1 : out std_logic;
	      ENA_2 : out std_logic);
    end component;
	--IP (Intellectual Property) of the RAM
	component blk_mem_gen_0 is
    PORT (
        clka : IN STD_LOGIC;
         ena : IN STD_LOGIC;
         wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
       addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
        dina : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        clkb : IN STD_LOGIC;
         enb : IN STD_LOGIC;
       addrb : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
       doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    end component;
	--Define the "wires" to join the components
	signal RESET_UART : std_logic;
	signal READY : std_logic;
	signal DATA : std_logic_vector(7 downto 0);
	signal ENA_1, ENA_2 : std_logic;
	signal ENB_1, ENB_2 : std_logic;
	signal ADDA, ADDB_1, ADDB_2 : std_logic_vector(9 downto 0);
	signal DOUTB_1, DOUTB_2 : std_logic_vector(7 downto 0);
	signal CV, CH : std_logic_vector(9 downto 0);
begin
    RESET_UART <= NOT RESET; --The UART DRIVER RESET is activated for 0 logic value
	--UART-RAM memory writer
	CONTROLLER_UART: CONTROL_UART port map(
	    READY => READY,
		RESET => RESET,
		  CLK => CLK,
		 DATA => DATA,
		 ADDA => ADDA,
		ENA_1 => ENA_1,
		ENA_2 => ENA_2);
	--UART DRIVER
	UART_DIVER: UART_RX port map(
	       reset => RESET_UART,
             clk => CLK,
		      rx => RX,
		data_out => DATA,
		   ready => READY);
	--Memory RAM Block 1
	RAM_1: blk_mem_gen_0 port map(
	     clka => CLK,
		 clkb => CLK,
		  ena => ENA_1,
		  wea(0) => ENA_1,
		addra => ADDA,
		 dina => DATA,
		  enb => ENB_1,
		addrb => ADDB_1,
		doutb => DOUTB_1);
	--Memory RAM Block 2
    RAM_2: blk_mem_gen_0 port map(
	     clka => CLK,
		 clkb => CLK,
		  ena => ENA_2,
		  wea(0) => ENA_2,
		addra => ADDA,
		 dina => DATA,
		  enb => ENB_2,
		addrb => ADDB_2,
		doutb => DOUTB_2);
	--Controller of the VGA
	CONTROLLER_VGA: CONTROL_VGA port map(
	      CLK => CLK,
		RESET => RESET,
		 CH_o => CH,
		 CV_o => CV,
		HSYNC => HSYNC,
		VSYNC => VSYNC);
	--Data Path to communicate the values written in the RAM memory with a VGA screen
	DATA_PATH_1: VGA_DATA port map(
	      CLK => CLK,
		RESET => RESET,
		   CH => CH,
		   CV => CV,
		 ADDB => ADDB_1,
		  ENB => ENB_1,
		DOUTB => DOUTB_1,
		COLOR => COLOR_R);
	DATA_PATH_2: VGA_DATA port map(
	      CLK => CLK,
		RESET => RESET,
		   CH => CH,
		   CV => CV,
		 ADDB => ADDB_2,
		  ENB => ENB_2,
		DOUTB => DOUTB_2,
		COLOR => COLOR_G);
	DATA_PATH_3: VGA_DATA port map(
	      CLK => CLK,
		RESET => RESET,
		   CH => CH,
		   CV => CV,
		--ADDB => ADDB_2,
		--ENB => ENB_2,
		DOUTB => "01111111", --Ground line printed
		COLOR => COLOR_B);
end A1;
